// Copyright (c) 2023 Conless Pan

// This source code is licensed under the MIT license found in the
// LICENSE file in the root directory of this source tree.

// This file contains the implementation of the fetch scheduler of the Gelato GPU. It chooses a warp in the pc table when the fetch unit is ready to fetch a new instruction.

`include "gelato_macros.svh"
`include "gelato_types.svh"

import gelato_types::*;

module gelato_fetch_scheduler (
  input logic clk,
  input logic rst_n,
  input logic rdy,

  // Get the pc of each warp
  gelato_pctable_fetchskd_if.slave pc_table_if,
  // Receive the buffer information
  gelato_ibuffer_fetchskd_if.slave ibuffer_if,

  // Send the pc to the fetch unit
  output logic dout_valid,
  input logic dout_ready,
  output pc_info_t dout
);
  //============================================================================
  // Information of each warp. delivered by the pc table and instruction buffer
  //============================================================================
  logic [`WARP_NUM-1:0] valid;
  logic [`WARP_NUM-1:0] warp_disabled;

  generate
    for (genvar i = 0; i < `WARP_NUM; i++) begin : gen_warp_valid
      assign valid[i] = pc_table_if.valid[i] && !warp_disabled[i] && ibuffer_if.available[i];
    end
  endgenerate

  always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      warp_disabled <= 0;
    end else if (pc_table_if.activate_valid) begin
      warp_disabled[pc_table_if.activate_warp_num] <= 0;
    end
  end

  //============================================================================
  // Selected warp number, generated by the round arbiter
  //============================================================================
  warp_num_t selected_warp;
  logic selected_valid;
  addr_t selected_pc;
  split_table_num_t selected_split_table_num;

  gelato_round_arbiter #(
    .PORT_NUM_WIDTH(`WARP_NUM_WIDTH),
    .STEP_LENGTH(2)
  ) round_arbiter (
    .clk(clk),
    .rst_n(rst_n),
    .req(valid),
    .selected(selected_warp)
  );

  assign selected_valid = valid[selected_warp];
  assign selected_pc = pc_table_if.pc[selected_warp];
  assign selected_split_table_num = pc_table_if.split_table_num[selected_warp];

  //============================================================================
  // Transition of state
  //============================================================================
  typedef enum logic { GENERATE_PC, WAIT_READY } state_t;
  state_t state_q, state_d;

  always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      state_q <= GENERATE_PC;
    end else begin
      state_q <= state_d;
    end
  end

  //============================================================================
  // Condition of state transition
  //============================================================================
  always_comb begin
    case (state_q)
      GENERATE_PC: begin
        state_d = selected_valid ? WAIT_READY : GENERATE_PC;
      end
      WAIT_READY: begin
        state_d = dout_ready ? GENERATE_PC : WAIT_READY;
      end
      default: begin
        $fatal(0, "gelato_fetch_scheduler: Invalid state");
      end
    endcase
  end

  //============================================================================
  // Output
  //============================================================================
  always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      dout_valid <= 0;
    end else begin
      case (state_d)
        GENERATE_PC: begin
          dout_valid <= 0;
        end
        WAIT_READY: begin
          dout_valid <= 1;
          dout.warp_num <= selected_warp;
          dout.pc <= selected_pc;
          dout.split_table_num <= selected_split_table_num;
        end
        default: begin
          $fatal(0, "gelato_fetch_scheduler: Invalid state");
        end
      endcase
    end
  end
endmodule
